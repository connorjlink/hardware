`include "../util/register.v"

module eauD_A(input[7:0] d, input di, clk, hs, ls, ao, output[15:0] a);

endmodule


module eau_A_D(input[15:0] a, input ai, clk, hs, ls, do, output[7:0] d);

endmodule