//decoder block
//this module is basically a wrapper on embedded microcode

module db
(
    input[7:0] insn, d1, d2, d3,

    input clk, rst,
);

    reg[31:0] ucode[255:0];

    initial 
    begin

    end

    always @()


endmodule