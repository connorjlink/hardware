//this module is basically a wrapper on embedded microcode

module db
(
    input[7:0] insn, d1, d2, d3
);

    reg[31:0] ucode[255:0];


endmodule