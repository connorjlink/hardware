`include "../util/mux/mux_8b.v"

module shift_8b(input[7:0] a, input[2:0] b, input lr, output[7:0] o);


endmodule