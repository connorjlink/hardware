module not_1b(input a, output b);
    assign b = ~a;
endmodule