module not_1w(input a, output b);
    assign b = ~a;
endmodule