module or_3w(input a, b, c, output d);
    assign d = (a | b | c);
endmodule