module mux_2b(input a, b, c, d, input[1:0] s, output o);

endmodule