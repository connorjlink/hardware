module cpu
(

);


endmodule