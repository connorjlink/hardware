module or_2w(input a, b, output c);
    assign c = (a | b);
endmodule