`timescale 1ns / 100ps
`include "lsu.v"

module lsu_tb;


endmodule