module and_2w(input a, b, output c);
    assign c = (a & b);
endmodule