module and_1b(input a, b, output c);
    assign c = (a & b);
endmodule